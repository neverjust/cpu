`timescale 1ns / 1ps
module CLA_4(X,Y,Cin,S,Cout);
    input [3:0]X,Y;
    input Cin;
    output [3:0]S;
    output Cout;
    or j0(J0,X[0],Y[0]);
    or j1(J1,X[1],Y[1]);
    or j2(J2,X[2],Y[2]);
    or j3(J3,X[3],Y[3]);
    and i0(I0,X[0],Y[0]);
    and i1(I1,X[1],Y[1]);
    and i2(I2,X[2],Y[2]);
    and i3(I3,X[3],Y[3]);
    not u0(U0,I0);
    not u1(U1,I1);
    not u2(U2,I2);
    not u3(U3,I3);
    and i4(I4,U0,J0);
    and i5(I5,U1,J1);
    and i6(I6,U2,J2);
    and i7(I7,U3,J3);
    nand v0(V0,Cin,J0);
    nand v1(V1,Cin,J0,J1);
    nand v2(V2,I0,J1);
    nand v3(V3,Cin,J0,J1,J2);
    nand v4(V4,I0,J1,J2);
    nand v5(V5,I1,J2);
    nand v6(V6,Cin,J0,J1,J2,J3);
    nand v7(V7,I0,J1,J2,J3);
    nand v8(V8,I1,J2,J3);
    nand v9(V9,I2,J3);
    nand v10(V10,V0,U0);
    nand v11(V11,V1,V2,U1);
    nand v12(V12,V3,V4,V5,U2);
    nand v13(Cout,V6,V7,V8,V9,U3);
    xor m0(S[0],Cin,I4);
    xor m1(S[1],V10,I5);
    xor m2(S[2],V11,I6);
    xor m3(S[3],V12,I7);
endmodule
